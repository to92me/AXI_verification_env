
package dut_testing_test_and_seqs_pkq;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "dut_testing/testing/sequences/dut_register_model_base_sequence.sv"


endpackage

`endif