module name;
	
endmodule
