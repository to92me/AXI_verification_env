//This is dummy DUT. 

module dut( input axi_clock, input axi_reset, axi_if axi_if);

endmodule