package name;
	
endpackage
