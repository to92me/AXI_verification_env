`ifndef DUT_TESTING_TYPES
`define DUT_TESTING_TYPES

typedef dut_testing_logger_results logger_result_queue[$];

`endif