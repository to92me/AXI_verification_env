
`ifndef TEST_PKG_SV
`define TEST_PKG_SV


//package test_pkg;
/*
	// ==================== SEQUENCES =============================
	typedef class dut_register_model_base_sequence;
	typedef class count_seq;
	typedef class dut_register_model_test_sequence;

	// ============================================================

	// ====================== TESTS ===============================
	typedef class dut_register_model_test_base;

	// ============================================================

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "axi_uvc/sv/axi_pkg.sv"
	import axi_pkg::*;

	`include "dut_register_layer/sv/dut_register_model_pkg.sv"
	import dut_register_model_pkg::*;

	`include "dut_testing/sv/register_model_env_pkg.sv"
	import register_model_env_pkg::*;

	// ==================== SEQUENCES =============================
	`include "dut_testing/testing/sequences/count_seq.sv"
	`include "dut_testing/testing/sequences/dut_register_model_base_sequence.sv"

	// ============================================================

	// ====================== TESTS ===============================
	`include "dut_testing/sv/test_tb/test.sv"

	// ============================================================
*/
//endpackage

`endif