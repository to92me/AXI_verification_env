`ifndef DUT_REGISTER_MODEL_TEST_PKG_SVH
`define DUT_REGISTER_MODEL_TEST_PKG_SVH

package uvc_company_uvc_name_pkg;


endpackage



`endif