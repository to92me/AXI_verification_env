/******************************************************************************
	* DVT CODE TEMPLATE: interface
	* Created by root on Aug 2, 2015
	* ovc_company = ovc_company, ovc_name = ovc_name ovc_if = ovc_if
	* interface arguments = interface_args
*******************************************************************************/

//-------------------------------------------------------------------------
//
// INTERFACE: ovc_company_ovc_name_ovc_if
//
//-------------------------------------------------------------------------

interface ovc_company_ovc_name_ovc_if (interface_args);

	// TODO: Define the interface signals here
	

endinterface : ovc_company_ovc_name_ovc_if
